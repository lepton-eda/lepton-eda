*
.model unknown_LVD (stuff)
