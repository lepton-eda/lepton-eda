LIBRARY ieee,disciplines;
USE ieee.math_real.all;
USE ieee.math_real.all;
USE work.electrical_system.all;
USE work.all;
-- Entity declaration -- 

ENTITY bjt_transistor_simple_top IS
END ENTITY bjt_transistor_simple_top; 

