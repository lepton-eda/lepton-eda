.model
D
