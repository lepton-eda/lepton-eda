;
; This file is really a gnetlistrc file.
; It is renamed to gnetlistrc before any vhdl backend test is run.
;
; The path is hardcoded for now.
;

(component-library "${HOME}/geda/share/gEDA/sym/vhdl")


